tb
`timescale 1ns / 1ps

module fft64pt_stage1_tb;

    // Testbench signals
    reg clk;
    reg signed [1:0] r[0:63];
    reg signed [1:0] i[0:63];
    wire signed [44:0] R[0:63];
    wire signed [44:0] I[0:63];

    // Instantiate the DUT (Device Under Test)
    fft64pt_stage1 dut (
        .clk(clk),
        .r0(r[0]), .r1(r[1]), .r2(r[2]), .r3(r[3]), .r4(r[4]), .r5(r[5]), .r6(r[6]), .r7(r[7]),
        .r8(r[8]), .r9(r[9]), .r10(r[10]), .r11(r[11]), .r12(r[12]), .r13(r[13]), .r14(r[14]), .r15(r[15]),
        .r16(r[16]), .r17(r[17]), .r18(r[18]), .r19(r[19]), .r20(r[20]), .r21(r[21]), .r22(r[22]), .r23(r[23]),
        .r24(r[24]), .r25(r[25]), .r26(r[26]), .r27(r[27]), .r28(r[28]), .r29(r[29]), .r30(r[30]), .r31(r[31]),
        .r32(r[32]), .r33(r[33]), .r34(r[34]), .r35(r[35]), .r36(r[36]), .r37(r[37]), .r38(r[38]), .r39(r[39]),
        .r40(r[40]), .r41(r[41]), .r42(r[42]), .r43(r[43]), .r44(r[44]), .r45(r[45]), .r46(r[46]), .r47(r[47]),
        .r48(r[48]), .r49(r[49]), .r50(r[50]), .r51(r[51]), .r52(r[52]), .r53(r[53]), .r54(r[54]), .r55(r[55]),
        .r56(r[56]), .r57(r[57]), .r58(r[58]), .r59(r[59]), .r60(r[60]), .r61(r[61]), .r62(r[62]), .r63(r[63]),
        .i0(i[0]), .i1(i[1]), .i2(i[2]), .i3(i[3]), .i4(i[4]), .i5(i[5]), .i6(i[6]), .i7(i[7]),
        .i8(i[8]), .i9(i[9]), .i10(i[10]), .i11(i[11]), .i12(i[12]), .i13(i[13]), .i14(i[14]), .i15(i[15]),
        .i16(i[16]), .i17(i[17]), .i18(i[18]), .i19(i[19]), .i20(i[20]), .i21(i[21]), .i22(i[22]), .i23(i[23]),
        .i24(i[24]), .i25(i[25]), .i26(i[26]), .i27(i[27]), .i28(i[28]), .i29(i[29]), .i30(i[30]), .i31(i[31]),
        .i32(i[32]), .i33(i[33]), .i34(i[34]), .i35(i[35]), .i36(i[36]), .i37(i[37]), .i38(i[38]), .i39(i[39]),
        .i40(i[40]), .i41(i[41]), .i42(i[42]), .i43(i[43]), .i44(i[44]), .i45(i[45]), .i46(i[46]), .i47(i[47]),
        .i48(i[48]), .i49(i[49]), .i50(i[50]), .i51(i[51]), .i52(i[52]), .i53(i[53]), .i54(i[54]), .i55(i[55]),
        .i56(i[56]), .i57(i[57]), .i58(i[58]), .i59(i[59]), .i60(i[60]), .i61(i[61]), .i62(i[62]), .i63(i[63]),
        .R0(R[0]), .R1(R[1]), .R2(R[2]), .R3(R[3]), .R4(R[4]), .R5(R[5]), .R6(R[6]), .R7(R[7]),
        .R8(R[8]), .R9(R[9]), .R10(R[10]), .R11(R[11]), .R12(R[12]), .R13(R[13]), .R14(R[14]), .R15(R[15]),
        .R16(R[16]), .R17(R[17]), .R18(R[18]), .R19(R[19]), .R20(R[20]), .R21(R[21]), .R22(R[22]), .R23(R[23]),
        .R24(R[24]), .R25(R[25]), .R26(R[26]), .R27(R[27]), .R28(R[28]), .R29(R[29]), .R30(R[30]), .R31(R[31]),
        .R32(R[32]), .R33(R[33]), .R34(R[34]), .R35(R[35]), .R36(R[36]), .R37(R[37]), .R38(R[38]), .R39(R[39]),
        .R40(R[40]), .R41(R[41]), .R42(R[42]), .R43(R[43]), .R44(R[44]), .R45(R[45]), .R46(R[46]), .R47(R[47]),
        .R48(R[48]), .R49(R[49]), .R50(R[50]), .R51(R[51]), .R52(R[52]), .R53(R[53]), .R54(R[54]), .R55(R[55]),
        .R56(R[56]), .R57(R[57]), .R58(R[58]), .R59(R[59]), .R60(R[60]), .R61(R[61]), .R62(R[62]), .R63(R[63]),
        .I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .I4(I[4]), .I5(I[5]), .I6(I[6]), .I7(I[7]),
        .I8(I[8]), .I9(I[9]), .I10(I[10]), .I11(I[11]), .I12(I[12]), .I13(I[13]), .I14(I[14]), .I15(I[15]),
        .I16(I[16]), .I17(I[17]), .I18(I[18]), .I19(I[19]), .I20(I[20]), .I21(I[21]), .I22(I[22]), .I23(I[23]),
        .I24(I[24]), .I25(I[25]), .I26(I[26]), .I27(I[27]), .I28(I[28]), .I29(I[29]), .I30(I[30]), .I31(I[31]),
        .I32(I[32]), .I33(I[33]), .I34(I[34]), .I35(I[35]), .I36(I[36]), .I37(I[37]), .I38(I[38]), .I39(I[39]),
        .I40(I[40]), .I41(I[41]), .I42(I[42]), .I43(I[43]), .I44(I[44]), .I45(I[45]), .I46(I[46]), .I47(I[47]),
        .I48(I[48]), .I49(I[49]), .I50(I[50]), .I51(I[51]), .I52(I[52]), .I53(I[53]), .I54(I[54]), .I55(I[55]),
        .I56(I[56]), .I57(I[57]), .I58(I[58]), .I59(I[59]), .I60(I[60]), .I61(I[61]), .I62(I[62]), .I63(I[63])
    );

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk;  // 10ns clock period
    end

    // Initialize input signals without using a loop
    initial begin
        // Manually set input values

    // Manually set input values for each element
    r[0] = 2'b00; i[0] = 2'b00;
    r[1] = 2'b01; i[1] = 2'b01;
    r[2] = 2'b10; i[2] = 2'b10;
    r[3] = 2'b11; i[3] = 2'b11;
    r[4] = 2'b00; i[4] = 2'b01;
    r[5] = 2'b01; i[5] = 2'b10;
    r[6] = 2'b10; i[6] = 2'b11;
    r[7] = 2'b11; i[7] = 2'b00;
    r[8] = 2'b00; i[8] = 2'b11;
    r[9] = 2'b01; i[9] = 2'b10;
    r[10] = 2'b10; i[10] = 2'b01;
    r[11] = 2'b11; i[11] = 2'b00;
    r[12] = 2'b00; i[12] = 2'b01;
    r[13] = 2'b01; i[13] = 2'b11;
    r[14] = 2'b10; i[14] = 2'b00;
    r[15] = 2'b11; i[15] = 2'b10;
    r[16] = 2'b00; i[16] = 2'b10;
    r[17] = 2'b01; i[17] = 2'b00;
    r[18] = 2'b10; i[18] = 2'b11;
    r[19] = 2'b11; i[19] = 2'b01;
    r[20] = 2'b00; i[20] = 2'b11;
    r[21] = 2'b01; i[21] = 2'b10;
    r[22] = 2'b10; i[22] = 2'b01;
    r[23] = 2'b11; i[23] = 2'b00;
    r[24] = 2'b00; i[24] = 2'b01;
    r[25] = 2'b01; i[25] = 2'b10;
    r[26] = 2'b10; i[26] = 2'b11;
    r[27] = 2'b11; i[27] = 2'b00;
    r[28] = 2'b00; i[28] = 2'b11;
    r[29] = 2'b01; i[29] = 2'b10;
    r[30] = 2'b10; i[30] = 2'b01;
    r[31] = 2'b11; i[31] = 2'b00;
    r[32] = 2'b00; i[32] = 2'b01;
    r[33] = 2'b01; i[33] = 2'b11;
    r[34] = 2'b10; i[34] = 2'b00;
    r[35] = 2'b11; i[35] = 2'b10;
    r[36] = 2'b00; i[36] = 2'b10;
    r[37] = 2'b01; i[37] = 2'b00;
    r[38] = 2'b10; i[38] = 2'b11;
    r[39] = 2'b11; i[39] = 2'b01;
    r[40] = 2'b00; i[40] = 2'b11;
    r[41] = 2'b01; i[41] = 2'b10;
    r[42] = 2'b10; i[42] = 2'b01;
    r[43] = 2'b11; i[43] = 2'b00;
    r[44] = 2'b00; i[44] = 2'b01;
    r[45] = 2'b01; i[45] = 2'b10;
    r[46] = 2'b10; i[46] = 2'b11;
    r[47] = 2'b11; i[47] = 2'b00;
    r[48] = 2'b00; i[48] = 2'b11;
    r[49] = 2'b01; i[49] = 2'b10;
    r[50] = 2'b10; i[50] = 2'b01;
    r[51] = 2'b11; i[51] = 2'b00;
    r[52] = 2'b00; i[52] = 2'b01;
    r[53] = 2'b01; i[53] = 2'b11;
    r[54] = 2'b10; i[54] = 2'b00;
    r[55] = 2'b11; i[55] = 2'b10;
    r[56] = 2'b00; i[56] = 2'b10;
    r[57] = 2'b01; i[57] = 2'b00;
    r[58] = 2'b10; i[58] = 2'b11;
    r[59] = 2'b11; i[59] = 2'b01;
    r[60] = 2'b00; i[60] = 2'b11;
    r[61] = 2'b01; i[61] = 2'b10;
    r[62] = 2'b10; i[62] = 2'b01;
    r[63] = 2'b11; i[63] = 2'b00;

    // Wait for some time to observe output

        // Observe for some cycles
        #1000 $stop;
    end

endmodule